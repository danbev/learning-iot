module first(input BUT1, output LED1);

  assign LED1 = BUT1;

endmodule
