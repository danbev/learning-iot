module first(input BUT1, LED1);
  assign LED1 = BUT1;
endmodule
